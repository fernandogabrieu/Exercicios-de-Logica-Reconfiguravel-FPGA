----------------------------------------------------
-- Código top-level calc.vhd
----------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.all;
LIBRARY work;
USE work.package_calculadora.all;


------------------------------------------------------------------------------------------------------------------------------------------------------------
ENTITY CALC IS
	PORT(A : IN INTEGER RANGE 0 TO 7;
		  B : IN INTEGER RANGE 0 TO 7;
		  SEL : IN std_logic;
		  OUTPUT : OUT INTEGER RANGE 0 TO 63); 
END CALC;

------------------------------------------------------------------------------------------------------------------------------------------------------------

ARCHITECTURE logic of CALC IS
BEGIN
	calculadora(A, B, SEL, OUTPUT);
END logic;
------------------------------------------------------------------------------------------------------------------------------------------------------------

